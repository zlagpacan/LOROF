/*
    Filename: bcb_wrapper.sv
    Author: zlagpacan
    Description: RTL wrapper around bcb module. 
    Spec: LOROF/spec/design/bcb.md
*/

`timescale 1ns/100ps

`include "corep.vh"

module bcb_wrapper #(
) (

    // seq
    input logic CLK,
    input logic nRST,


    // save control
	input logic next_save_valid,
	input corep::bcb_info_t next_save_bcb_info,

	output corep::bcb_idx_t last_save_bcb_idx,

    // restore control
	input corep::bcb_idx_t next_restore_bcb_idx,

	output corep::bcb_info_t last_restore_bcb_info
);

    // ----------------------------------------------------------------
    // Direct Module Connections:


    // save control
	logic save_valid;
	corep::bcb_info_t save_bcb_info;

	corep::bcb_idx_t save_bcb_idx;

    // restore control
	corep::bcb_idx_t restore_bcb_idx;

	corep::bcb_info_t restore_bcb_info;

    // ----------------------------------------------------------------
    // Module Instantiation:

	bcb #(
	) WRAPPED_MODULE (.*);

    // ----------------------------------------------------------------
    // Wrapper Registers:

    always_ff @ (posedge CLK, negedge nRST) begin
        if (~nRST) begin


		    // save control
			save_valid <= '0;
			save_bcb_info <= '0;

			last_save_bcb_idx <= '0;

		    // restore control
			restore_bcb_idx <= '0;

			last_restore_bcb_info <= '0;
        end
        else begin


		    // save control
			save_valid <= next_save_valid;
			save_bcb_info <= next_save_bcb_info;

			last_save_bcb_idx <= save_bcb_idx;

		    // restore control
			restore_bcb_idx <= next_restore_bcb_idx;

			last_restore_bcb_info <= restore_bcb_info;
        end
    end

endmodule