/*
    Filename: instr_types.vh
    Author: zlagpacan
    Description: Package Header File for Instruction Types
*/

`ifndef INSTR_TYPES_VH
`define INSTR_TYPES_VH

package instr_types;

    // ----------------------------------------------------------------
    // Custom op decoding:

    // TODO: finish op encoding in instr_list.md

endpackage

`endif // CORE_TYPES_VH