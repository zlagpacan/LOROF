// need to send decode_unit restart to fetch_unit AFTER decode_unit update has finished
    // don't want another mispred