/*
    Filename: alu_iq_tb.sv
    Author: zlagpacan
    Description: Testbench for alu_iq module. 
    Spec: LOROF/spec/design/alu_iq.md
*/

`timescale 1ns/100ps

`include "core_types_pkg.vh"
import core_types_pkg::*;

module alu_iq_tb ();

    ///////////////////////////////////////////////////////////////////////////////////////////////////////
    // TB setup:

    // parameters
    parameter PERIOD = 10;

    // TB signals:
    logic CLK = 1'b1, nRST;
    string test_case;
    string sub_test_case;
    int test_num = 0;
    int num_errors = 0;
    logic tb_error = 1'b0;

    // clock gen
    always begin #(PERIOD/2); CLK = ~CLK; end

    ///////////////////////////////////////////////////////////////////////////////////////////////////////
    // DUT signals:


    // ALU op dispatch by entry
	logic [3:0] tb_dispatch_valid_by_entry;
	logic [3:0][3:0] tb_dispatch_op_by_entry;
	logic [3:0][31:0] tb_dispatch_imm_by_entry;
	logic [3:0][LOG_PR_COUNT-1:0] tb_dispatch_A_PR_by_entry;
	logic [3:0] tb_dispatch_A_unneeded_by_entry;
	logic [3:0] tb_dispatch_A_ready_by_entry;
	logic [3:0][LOG_PR_COUNT-1:0] tb_dispatch_B_PR_by_entry;
	logic [3:0] tb_dispatch_is_imm_by_entry;
	logic [3:0] tb_dispatch_B_ready_by_entry;
	logic [3:0][LOG_PR_COUNT-1:0] tb_dispatch_dest_PR_by_entry;

    // ALU op dispatch feedback by entry
    logic [3:0] DUT_dispatch_open_by_entry, expected_dispatch_open_by_entry;

    // ALU pipeline feedback
    logic tb_pipeline_ready;

    // writeback bus
	logic [PRF_BANK_COUNT-1:0] tb_WB_valid_by_bank;
	logic [PRF_BANK_COUNT-1:0][LOG_PR_COUNT-LOG_PRF_BANK_COUNT-1:0] tb_WB_upper_PR_by_bank;

    // ALU op issue to ALU pipeline
	logic DUT_issue_valid, expected_issue_valid;
	logic [3:0] DUT_issue_op, expected_issue_op;
	logic DUT_issue_is_imm, expected_issue_is_imm;
	logic [31:0] DUT_issue_imm, expected_issue_imm;
	logic DUT_issue_A_unneeded, expected_issue_A_unneeded;
	logic DUT_issue_A_forward, expected_issue_A_forward;
	logic [LOG_PRF_BANK_COUNT-1:0] DUT_issue_A_bank, expected_issue_A_bank;
	logic DUT_issue_B_forward, expected_issue_B_forward;
	logic [LOG_PRF_BANK_COUNT-1:0] DUT_issue_B_bank, expected_issue_B_bank;
	logic [LOG_PR_COUNT-1:0] DUT_issue_dest_PR, expected_issue_dest_PR;

    // reg read req to PRF
	logic DUT_PRF_req_A_valid, expected_PRF_req_A_valid;
	logic [LOG_PR_COUNT-1:0] DUT_PRF_req_A_PR, expected_PRF_req_A_PR;
	logic DUT_PRF_req_B_valid, expected_PRF_req_B_valid;
	logic [LOG_PR_COUNT-1:0] DUT_PRF_req_B_PR, expected_PRF_req_B_PR;

    ///////////////////////////////////////////////////////////////////////////////////////////////////////
    // DUT instantiation:

	alu_iq DUT (

		// seq
		.CLK(CLK),
		.nRST(nRST),

	    // ALU op dispatch by entry
		.dispatch_valid_by_entry(tb_dispatch_valid_by_entry),
		.dispatch_op_by_entry(tb_dispatch_op_by_entry),
		.dispatch_imm_by_entry(tb_dispatch_imm_by_entry),
		.dispatch_A_PR_by_entry(tb_dispatch_A_PR_by_entry),
		.dispatch_A_unneeded_by_entry(tb_dispatch_A_unneeded_by_entry),
		.dispatch_A_ready_by_entry(tb_dispatch_A_ready_by_entry),
		.dispatch_B_PR_by_entry(tb_dispatch_B_PR_by_entry),
		.dispatch_is_imm_by_entry(tb_dispatch_is_imm_by_entry),
		.dispatch_B_ready_by_entry(tb_dispatch_B_ready_by_entry),
		.dispatch_dest_PR_by_entry(tb_dispatch_dest_PR_by_entry),

        // ALU op dispatch feedback by entry
        .dispatch_open_by_entry(DUT_dispatch_open_by_entry),

        // ALU pipeline feedback
        .pipeline_ready(tb_pipeline_ready),

	    // writeback bus
		.WB_valid_by_bank(tb_WB_valid_by_bank),
		.WB_upper_PR_by_bank(tb_WB_upper_PR_by_bank),

	    // ALU op issue to ALU pipeline
		.issue_valid(DUT_issue_valid),
		.issue_op(DUT_issue_op),
		.issue_is_imm(DUT_issue_is_imm),
		.issue_imm(DUT_issue_imm),
		.issue_A_unneeded(DUT_issue_A_unneeded),
		.issue_A_forward(DUT_issue_A_forward),
		.issue_A_bank(DUT_issue_A_bank),
		.issue_B_forward(DUT_issue_B_forward),
		.issue_B_bank(DUT_issue_B_bank),
		.issue_dest_PR(DUT_issue_dest_PR),

	    // reg read req to PRF
		.PRF_req_A_valid(DUT_PRF_req_A_valid),
		.PRF_req_A_PR(DUT_PRF_req_A_PR),
		.PRF_req_B_valid(DUT_PRF_req_B_valid),
		.PRF_req_B_PR(DUT_PRF_req_B_PR)
	);

    ///////////////////////////////////////////////////////////////////////////////////////////////////////
    // tasks:

    task check_outputs();
    begin
		if (expected_dispatch_open_by_entry !== DUT_dispatch_open_by_entry) begin
			$display("TB ERROR: expected_dispatch_open_by_entry (%h) != DUT_dispatch_open_by_entry (%h)",
				expected_dispatch_open_by_entry, DUT_dispatch_open_by_entry);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_valid !== DUT_issue_valid) begin
			$display("TB ERROR: expected_issue_valid (%h) != DUT_issue_valid (%h)",
				expected_issue_valid, DUT_issue_valid);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_op !== DUT_issue_op) begin
			$display("TB ERROR: expected_issue_op (%h) != DUT_issue_op (%h)",
				expected_issue_op, DUT_issue_op);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_is_imm !== DUT_issue_is_imm) begin
			$display("TB ERROR: expected_issue_is_imm (%h) != DUT_issue_is_imm (%h)",
				expected_issue_is_imm, DUT_issue_is_imm);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_imm !== DUT_issue_imm) begin
			$display("TB ERROR: expected_issue_imm (%h) != DUT_issue_imm (%h)",
				expected_issue_imm, DUT_issue_imm);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_A_unneeded !== DUT_issue_A_unneeded) begin
			$display("TB ERROR: expected_issue_A_unneeded (%h) != DUT_issue_A_unneeded (%h)",
				expected_issue_A_unneeded, DUT_issue_A_unneeded);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_A_forward !== DUT_issue_A_forward) begin
			$display("TB ERROR: expected_issue_A_forward (%h) != DUT_issue_A_forward (%h)",
				expected_issue_A_forward, DUT_issue_A_forward);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_A_bank !== DUT_issue_A_bank) begin
			$display("TB ERROR: expected_issue_A_bank (%h) != DUT_issue_A_bank (%h)",
				expected_issue_A_bank, DUT_issue_A_bank);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_B_forward !== DUT_issue_B_forward) begin
			$display("TB ERROR: expected_issue_B_forward (%h) != DUT_issue_B_forward (%h)",
				expected_issue_B_forward, DUT_issue_B_forward);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_B_bank !== DUT_issue_B_bank) begin
			$display("TB ERROR: expected_issue_B_bank (%h) != DUT_issue_B_bank (%h)",
				expected_issue_B_bank, DUT_issue_B_bank);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_issue_dest_PR !== DUT_issue_dest_PR) begin
			$display("TB ERROR: expected_issue_dest_PR (%h) != DUT_issue_dest_PR (%h)",
				expected_issue_dest_PR, DUT_issue_dest_PR);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_PRF_req_A_valid !== DUT_PRF_req_A_valid) begin
			$display("TB ERROR: expected_PRF_req_A_valid (%h) != DUT_PRF_req_A_valid (%h)",
				expected_PRF_req_A_valid, DUT_PRF_req_A_valid);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_PRF_req_A_PR !== DUT_PRF_req_A_PR) begin
			$display("TB ERROR: expected_PRF_req_A_PR (%h) != DUT_PRF_req_A_PR (%h)",
				expected_PRF_req_A_PR, DUT_PRF_req_A_PR);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_PRF_req_B_valid !== DUT_PRF_req_B_valid) begin
			$display("TB ERROR: expected_PRF_req_B_valid (%h) != DUT_PRF_req_B_valid (%h)",
				expected_PRF_req_B_valid, DUT_PRF_req_B_valid);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_PRF_req_B_PR !== DUT_PRF_req_B_PR) begin
			$display("TB ERROR: expected_PRF_req_B_PR (%h) != DUT_PRF_req_B_PR (%h)",
				expected_PRF_req_B_PR, DUT_PRF_req_B_PR);
			num_errors++;
			tb_error = 1'b1;
		end

        #(PERIOD / 10);
        tb_error = 1'b0;
    end
    endtask

    ///////////////////////////////////////////////////////////////////////////////////////////////////////
    // initial block:

    initial begin

        ///////////////////////////////////////////////////////////////////////////////////////////////////
        // reset:
        test_case = "reset";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

        // inputs:
        sub_test_case = "assert reset";
        $display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b0;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(posedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h0;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h0;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

        // inputs:
        sub_test_case = "deassert reset";
        $display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(posedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h0;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h0;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

        ///////////////////////////////////////////////////////////////////////////////////////////////////
        // simple chain:
        test_case = "simple chain";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: NOP", "\n\t\t",
            "dispatch2: NOP", "\n\t\t",
            "dispatch1: NOP", "\n\t\t",
            "dispatch0: ADD p3, p1:r, p2:r", "\n\t\t",
            "IQ3: NOP", "\n\t\t",
            "IQ2: NOP", "\n\t\t",
            "IQ1: NOP", "\n\t\t",
            "IQ0: NOP", "\n\t\t",
            "issue: NOP", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0001;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h1};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0001;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h2};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0001;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h3};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h0;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h0;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: NOP", "\n\t\t",
            "dispatch2: NOP", "\n\t\t",
            "dispatch1: NOP", "\n\t\t",
            "dispatch0: SLL p6, p4:f, p5:r", "\n\t\t",
            "IQ3: NOP", "\n\t\t",
            "IQ2: NOP", "\n\t\t",
            "IQ1: NOP", "\n\t\t",
            "IQ0: ADD p3, p1:r, p2:r", "\n\t\t",
            "issue: ADD p3, p1:r, p2:r", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0001;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0001};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h4};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h5};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0001;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h6};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h1;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h2;
		expected_issue_dest_PR = 6'h3;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b1;
		expected_PRF_req_A_PR = 6'h1;
		expected_PRF_req_B_valid = 1'b1;
		expected_PRF_req_B_PR = 6'h2;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: OR p12, p11:r, p8:f", "\n\t\t",
            "dispatch2: XORI p10, p8:f, 0xFFFFFFFF", "\n\t\t",
            "dispatch1: SLTI p9, p8:f, 0x678", "\n\t\t",
            "dispatch0: LUI p7, 0x12345000", "\n\t\t",
            "IQ3: NOP", "\n\t\t",
            "IQ2: NOP", "\n\t\t",
            "IQ1: NOP", "\n\t\t",
            "IQ0: v SLL p6, p4:F, p5:r", "\n\t\t",
            "issue: SLL p6, p4:F, p5:r", "\n\t\t",
			"activity: WB p4", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b1111;
		tb_dispatch_op_by_entry = {4'b0110, 4'b0100, 4'b0010, 4'b1111};
		tb_dispatch_imm_by_entry = {32'h0, 32'hFFFFFFFF, 32'h678, 32'h12345000};
		tb_dispatch_A_PR_by_entry = {6'hB, 6'h8, 6'h8, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0001;
		tb_dispatch_A_ready_by_entry = 4'b1000;
		tb_dispatch_B_PR_by_entry = {6'h8, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0111;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'hC, 6'hA, 6'h9, 6'h7};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0001;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h1};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0001;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b1;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h1;
		expected_issue_dest_PR = 6'h6;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h4;
		expected_PRF_req_B_valid = 1'b1;
		expected_PRF_req_B_PR = 6'h5;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: v OR p12, p11:r, p8:f", "\n\t\t",
            "IQ2: v XORI p10, p8:f, 0xFFFFFFFF", "\n\t\t",
            "IQ1: v SLTI p9, p8:f, 0x678", "\n\t\t",
            "IQ0: v LUI p7, 0x12345000", "\n\t\t",
            "issue: i LUI p7, 0x12345000", "\n\t\t",
			"activity: pipeline not ready", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b0;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b0000;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b1111;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'h12345000;
		expected_issue_A_unneeded = 1'b1;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h7;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h0;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: v SRAI p14, p13:r, 0x123", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: v OR p12, p11:r, p8:f", "\n\t\t",
            "IQ2: v XORI p10, p8:f, 0xFFFFFFFF", "\n\t\t",
            "IQ1: v SLTI p9, p8:f, 0x678", "\n\t\t",
            "IQ0: v LUI p7, 0x12345000", "\n\t\t",
            "issue: v LUI p7, 0x12345000", "\n\t\t",
			"activity: ", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b1000;
		tb_dispatch_op_by_entry = {4'b1101, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h123, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'hD, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b1000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b1000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'hE, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1000;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b1111;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'h12345000;
		expected_issue_A_unneeded = 1'b1;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h7;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h0;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: v SRAI p14, p13:r, 0x123", "\n\t\t",
            "IQ2: v OR p12, p11:r, p8:f", "\n\t\t",
            "IQ1: v XORI p10, p8:f, 0xFFFFFFFF", "\n\t\t",
            "IQ0: v SLTI p9, p8:f, 0x678", "\n\t\t",
            "issue: v SRAI p14, p13:r, 0x123", "\n\t\t",
			"activity: ", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1000;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b1101;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'h123;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h1;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'hE;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b1;
		expected_PRF_req_A_PR = 6'hD;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: v OR p12, p11:r, p8:Fr", "\n\t\t",
            "IQ1: v XORI p10, p8:Fr, 0xFFFFFFFF", "\n\t\t",
            "IQ0: v SLTI p9, p8:F, 0x678", "\n\t\t",
            "issue: v SLTI p9, p8:F, 0x678", "\n\t\t",
			"activity: WB p8", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0001;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h2};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1100;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0010;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'h678;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b1;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h9;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h8;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: v SLTIU p19, p18:f, 0x543", "\n\t\t",
            "dispatch2: v OR p17, p15:f, p16:f", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: v OR p12, p11:r, p8:r", "\n\t\t",
            "IQ0: v XORI p10, p8:r, 0xFFFFFFFF", "\n\t\t",
            "issue: i XORI p10, p8:r, 0xFFFFFFFF", "\n\t\t",
			"activity: pipeline not ready", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b1100;
		tb_dispatch_op_by_entry = {4'b0011, 4'b0110, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h543, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h12, 6'hF, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h10, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b1000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h13, 6'h11, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b0;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1100;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0100;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'hFFFFFFFF;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'hA;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h8;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: v SLTIU p19, p18:f, 0x543", "\n\t\t",
            "IQ2: v OR p17, p15:f, p16:f", "\n\t\t",
            "IQ1: v OR p12, p11:r, p8:r", "\n\t\t",
            "IQ0: v XORI p10, p8:r, 0xFFFFFFFF", "\n\t\t",
            "issue: v XORI p10, p8:r, 0xFFFFFFFF", "\n\t\t",
			"activity: ", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0110, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1000;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0100;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'hFFFFFFFF;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'hA;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b1;
		expected_PRF_req_A_PR = 6'h8;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: v SLTIU p19, p18:f, 0x543", "\n\t\t",
            "IQ1: v OR p17, p15:f, p16:f", "\n\t\t",
            "IQ0: v OR p12, p11:r, p8:r", "\n\t\t",
            "issue: v OR p12, p11:r, p8:r", "\n\t\t",
			"activity: ", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0110, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1100;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0110;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h3;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'hC;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b1;
		expected_PRF_req_A_PR = 6'hB;
		expected_PRF_req_B_valid = 1'b1;
		expected_PRF_req_B_PR = 6'h8;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: v SLTIU p19, p18:Fr, 0x543", "\n\t\t",
            "IQ0: v OR p17, p15:F, p16:F", "\n\t\t",
            "issue: v OR p17, p15:F, p16:F", "\n\t\t",
			"activity: WB p15, p16, p18", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0110, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b1101;
		tb_WB_upper_PR_by_bank = {4'h3, 4'h4, 4'h0, 4'h4};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1110;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0110;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b1;
		expected_issue_A_bank = 2'h3;
		expected_issue_B_forward = 1'b1;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h11;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'hF;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h10;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: v ADD p27, p26:f, p26:f", "\n\t\t",
            "dispatch1: v SRL p25, p23:f, p24:f", "\n\t\t",
            "dispatch0: v SUB p22, p20:f, p21:f", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: i NOP", "\n\t\t",
            "IQ0: v SLTIU p19, p18:r, 0x543", "\n\t\t",
            "issue: v SLTIU p19, p18:r, 0x543", "\n\t\t",
			"activity: ", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0111;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0101, 4'b1000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h1A, 6'h17, 6'h14};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h1A, 6'h18, 6'h15};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h1B, 6'h19, 6'h16};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0011;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'h543;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h2;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h13;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b1;
		expected_PRF_req_A_PR = 6'h12;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: v ADD p27, p26:f, p26:f", "\n\t\t",
            "IQ1: v SRL p25, p23:f, p24:f", "\n\t\t",
            "IQ0: v SUB p22, p20:F, p21:F", "\n\t\t",
            "issue: v SUB p22, p20:F, p21:F", "\n\t\t",
			"activity: WB p20, p21", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0011;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h5, 4'h5};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1100;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b1000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b1;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b1;
		expected_issue_B_bank = 2'h1;
		expected_issue_dest_PR = 6'h16;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h14;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h15;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: v ADD p27, p26:f, p26:f", "\n\t\t",
            "IQ0: v SRL p25, p23:f, p24:Fr", "\n\t\t",
            "issue: i SRL p25, p23:f, p24:Fr", "\n\t\t",
			"activity: WB p24", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0001;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h6};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1100;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0101;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h3;
		expected_issue_B_forward = 1'b1;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h19;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h17;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h18;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: v ADD p27, p26:f, p26:f", "\n\t\t",
            "IQ0: v SRL p25, p23:F, p24:r", "\n\t\t",
            "issue: v SRL p25, p23:F, p24:r", "\n\t\t",
			"activity: WB p23", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b1000;
		tb_WB_upper_PR_by_bank = {4'h5, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1110;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0101;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b1;
		expected_issue_A_bank = 2'h3;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h19;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h17;
		expected_PRF_req_B_valid = 1'b1;
		expected_PRF_req_B_PR = 6'h18;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: i NOP", "\n\t\t",
            "IQ0: v ADD p27, p26:f, p26:f", "\n\t\t",
            "issue: i ADD p27, p26:f, p26:f", "\n\t\t",
			"activity: inv WB p26", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b1011;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h6, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1110;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h2;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h2;
		expected_issue_dest_PR = 6'h1B;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h1A;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h1A;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: v SLLI p29, p28:f, 0x3", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: i NOP", "\n\t\t",
            "IQ0: v ADD p27, p26:f, p26:f", "\n\t\t",
            "issue: v ADD p27, p26:f, p26:f", "\n\t\t",
			"activity: WB p26", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0001;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0001};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h3};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h1C};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0001;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h1D};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0100;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h6, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b1;
		expected_issue_A_bank = 2'h2;
		expected_issue_B_forward = 1'b1;
		expected_issue_B_bank = 2'h2;
		expected_issue_dest_PR = 6'h1B;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h1A;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h1A;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: i NOP", "\n\t\t",
            "IQ0: v SLLI p29, p28:Fr, 0x3", "\n\t\t",
            "issue: i SLLI p29, p28:Fr, 0x3", "\n\t\t",
			"activity: WB p28, pipeline not ready", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b0;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0001;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h7};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1110;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0001;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'h3;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b1;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h1D;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h1C;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: i NOP", "\n\t\t",
            "IQ0: v SLLI p29, p28:r, 0x3", "\n\t\t",
            "issue: v SLLI p29, p28:r, 0x3", "\n\t\t",
			"activity: ", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b1;
		expected_issue_op = 4'b0001;
		expected_issue_is_imm = 1'b1;
		expected_issue_imm = 32'h3;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h1D;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b1;
		expected_PRF_req_A_PR = 6'h1C;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

		@(posedge CLK);

		// inputs
		sub_test_case = {"\n\t\t", 
            "dispatch3: i NOP", "\n\t\t",
            "dispatch2: i NOP", "\n\t\t",
            "dispatch1: i NOP", "\n\t\t",
            "dispatch0: i NOP", "\n\t\t",
            "IQ3: i NOP", "\n\t\t",
            "IQ2: i NOP", "\n\t\t",
            "IQ1: i NOP", "\n\t\t",
            "IQ0: i NOP", "\n\t\t",
            "issue: i NOP", "\n\t\t",
			"activity: ", "\n\t\t"
        };
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // ALU op dispatch by entry
		tb_dispatch_valid_by_entry = 4'b0000;
		tb_dispatch_op_by_entry = {4'b0000, 4'b0000, 4'b0000, 4'b0000};
		tb_dispatch_imm_by_entry = {32'h0, 32'h0, 32'h0, 32'h0};
		tb_dispatch_A_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_A_unneeded_by_entry = 4'b0000;
		tb_dispatch_A_ready_by_entry = 4'b0000;
		tb_dispatch_B_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
		tb_dispatch_is_imm_by_entry = 4'b0000;
		tb_dispatch_B_ready_by_entry = 4'b0000;
		tb_dispatch_dest_PR_by_entry = {6'h0, 6'h0, 6'h0, 6'h0};
        // ALU op dispatch feedback by entry
        // ALU pipeline feedback
        tb_pipeline_ready = 1'b1;
	    // writeback bus
		tb_WB_valid_by_bank = 4'b0000;
		tb_WB_upper_PR_by_bank = {4'h0, 4'h0, 4'h0, 4'h0};
	    // ALU op issue to ALU pipeline
	    // reg read req to PRF

		@(negedge CLK);

		// outputs:

	    // ALU op dispatch by entry
        // ALU op dispatch feedback by entry
        expected_dispatch_open_by_entry = 4'b1111;
        // ALU pipeline feedback
	    // writeback bus
	    // ALU op issue to ALU pipeline
		expected_issue_valid = 1'b0;
		expected_issue_op = 4'b0000;
		expected_issue_is_imm = 1'b0;
		expected_issue_imm = 32'h0;
		expected_issue_A_unneeded = 1'b0;
		expected_issue_A_forward = 1'b0;
		expected_issue_A_bank = 2'h0;
		expected_issue_B_forward = 1'b0;
		expected_issue_B_bank = 2'h0;
		expected_issue_dest_PR = 6'h0;
	    // reg read req to PRF
		expected_PRF_req_A_valid = 1'b0;
		expected_PRF_req_A_PR = 6'h0;
		expected_PRF_req_B_valid = 1'b0;
		expected_PRF_req_B_PR = 6'h0;

		check_outputs();

        ///////////////////////////////////////////////////////////////////////////////////////////////////
        // finish:
        @(posedge CLK);
        
        test_case = "finish";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

        @(posedge CLK);

        $display();
        if (num_errors) begin
            $display("FAIL: %d tests fail", num_errors);
        end
        else begin
            $display("SUCCESS: all tests pass");
        end
        $display();

        $finish();
    end

endmodule

