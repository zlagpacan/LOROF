/*
  Module        : alu_pipeline
  UMV Component : System Verilog Assertions
  Author        : Adam Keith
*/

`ifndef ALU_PIPELINE_RST_SVA_SV
`define ALU_PIPELINE_RST_SVA_SV

// TODO:

`endif