/*
    Filename: bru_pred_info_updater_tb.sv
    Author: zlagpacan
    Description: Testbench for bru_pred_info_updater module. 
    Spec: LOROF/spec/design/bru_pred_info_updater.md
*/

`timescale 1ns/100ps

`include "core_types_pkg.vh"
import core_types_pkg::*;

module bru_pred_info_updater_tb ();

    // ----------------------------------------------------------------
    // TB setup:

    // parameters
    parameter PERIOD = 10;

    // TB signals:
    logic CLK = 1'b1, nRST;
    string test_case;
    string sub_test_case;
    int test_num = 0;
    int num_errors = 0;
    logic tb_error = 1'b0;

    // clock gen
    always begin #(PERIOD/2); CLK = ~CLK; end

    // ----------------------------------------------------------------
    // DUT signals:

    // inputs
	logic [3:0] tb_op;
	logic [BTB_PRED_INFO_WIDTH-1:0] tb_start_pred_info;
	logic tb_is_link_ra;
	logic tb_is_ret_ra;
	logic tb_is_taken;
	logic tb_is_mispredict;
	logic tb_is_out_of_range;

    // outputs
	logic [BTB_PRED_INFO_WIDTH-1:0] DUT_updated_pred_info, expected_updated_pred_info;

    // ----------------------------------------------------------------
    // DUT instantiation:

	bru_pred_info_updater DUT (

	    // inputs
		.op(tb_op),
		.start_pred_info(tb_start_pred_info),
		.is_link_ra(tb_is_link_ra),
		.is_ret_ra(tb_is_ret_ra),
		.is_taken(tb_is_taken),
		.is_mispredict(tb_is_mispredict),
		.is_out_of_range(tb_is_out_of_range),

	    // outputs
		.updated_pred_info(DUT_updated_pred_info)
	);

    // ----------------------------------------------------------------
    // tasks:

    task check_outputs();
    begin
		if (expected_updated_pred_info !== DUT_updated_pred_info) begin
			$display("TB ERROR: expected_updated_pred_info (%h) != DUT_updated_pred_info (%h)",
				expected_updated_pred_info, DUT_updated_pred_info);
			num_errors++;
			tb_error = 1'b1;
		end

        #(PERIOD / 10);
        tb_error = 1'b0;
    end
    endtask

    // ----------------------------------------------------------------
    // initial block:

    initial begin

        // ------------------------------------------------------------
        // reset:
        test_case = "reset";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

        // inputs:
        sub_test_case = "assert reset";
        $display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b0;
	    // inputs
		tb_op = 4'b0000;
		tb_start_pred_info = 8'h0;
		tb_is_link_ra = 1'b0;
		tb_is_ret_ra = 1'b0;
		tb_is_taken = 1'b0;
		tb_is_mispredict = 1'b0;
		tb_is_out_of_range = 1'b0;
	    // outputs

		@(posedge CLK); #(PERIOD/10);

		// outputs:

	    // inputs
	    // outputs
		expected_updated_pred_info = 8'b01000000;

		check_outputs();

        // inputs:
        sub_test_case = "deassert reset";
        $display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // inputs
		tb_op = 4'b0000;
		tb_start_pred_info = 8'h0;
		tb_is_link_ra = 1'b0;
		tb_is_ret_ra = 1'b0;
		tb_is_taken = 1'b0;
		tb_is_mispredict = 1'b0;
		tb_is_out_of_range = 1'b0;
	    // outputs

		@(posedge CLK); #(PERIOD/10);

		// outputs:

	    // inputs
	    // outputs
		expected_updated_pred_info = 8'b01000000;

		check_outputs();

        // ------------------------------------------------------------
        // basic coverage:
        test_case = "basic coverage";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "JALR !, 0(!) -> Jump";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // inputs
		tb_op = 4'b0000;
		tb_start_pred_info = 8'h0;
		tb_is_link_ra = 1'b0;
		tb_is_ret_ra = 1'b0;
		tb_is_taken = 1'b0;
		tb_is_mispredict = 1'b0;
		tb_is_out_of_range = 1'b0;
	    // outputs

		@(negedge CLK);

		// outputs:

	    // inputs
	    // outputs
		expected_updated_pred_info = 8'b01000000;

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "JALR ra, 0(!) -> JAL PC+4";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // inputs
		tb_op = 4'b0000;
		tb_start_pred_info = 8'h0;
		tb_is_link_ra = 1'b1;
		tb_is_ret_ra = 1'b0;
		tb_is_taken = 1'b0;
		tb_is_mispredict = 1'b0;
		tb_is_out_of_range = 1'b0;
	    // outputs

		@(negedge CLK);

		// outputs:

	    // inputs
	    // outputs
		expected_updated_pred_info = 8'b01011000;

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "JALR !, 0(ra) -> RET";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // inputs
		tb_op = 4'b0000;
		tb_start_pred_info = 8'h0;
		tb_is_link_ra = 1'b0;
		tb_is_ret_ra = 1'b1;
		tb_is_taken = 1'b0;
		tb_is_mispredict = 1'b0;
		tb_is_out_of_range = 1'b0;
	    // outputs

		@(negedge CLK);

		// outputs:

	    // inputs
	    // outputs
		expected_updated_pred_info = 8'b01100000;

		check_outputs();

        // ------------------------------------------------------------
        // finish:
        @(posedge CLK); #(PERIOD/10);
        
        test_case = "finish";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

        @(posedge CLK); #(PERIOD/10);

        $display();
        if (num_errors) begin
            $display("FAIL: %d tests fail", num_errors);
        end
        else begin
            $display("SUCCESS: all tests pass");
        end
        $display();

        $finish();
    end

endmodule