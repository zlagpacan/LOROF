// mq enq race condition: all mq entries younger than old mq entry trying to enq now
    // can keep timer in mq checking for too many cycles where
    // input enq ROB index older than all mq ROB index's