/*
    Filename: ras_tb.sv
    Author: zlagpacan
    Description: Testbench for ras module. 
    Spec: LOROF/spec/design/ras.md
*/

`timescale 1ns/100ps

`include "corep.vh"

module ras_tb #(
) ();

    // ----------------------------------------------------------------
    // TB setup:

    // parameters
    parameter PERIOD = 10;

    // TB signals:
    logic CLK = 1'b1, nRST;
    string test_case;
    string sub_test_case;
    int test_num = 0;
    int num_errors = 0;
    logic tb_error = 1'b0;

    // clock gen
    always begin #(PERIOD/2); CLK = ~CLK; end

    // ----------------------------------------------------------------
    // DUT signals:


    // pc_gen link control
	logic tb_link_valid;
	corep::PC38_t tb_link_pc38;

    // pc_gen return control
	logic tb_ret_valid;
	corep::PC38_t DUT_ret_pc38, expected_ret_pc38;
	corep::RAS_idx_t DUT_ret_ras_index, expected_ret_ras_index;

    // update control
	logic tb_update_valid;
	corep::RAS_idx_t tb_update_ras_index;

    // ----------------------------------------------------------------
    // DUT instantiation:

	ras #(
	) DUT (
		// seq
		.CLK(CLK),
		.nRST(nRST),


	    // pc_gen link control
		.link_valid(tb_link_valid),
		.link_pc38(tb_link_pc38),

	    // pc_gen return control
		.ret_valid(tb_ret_valid),
		.ret_pc38(DUT_ret_pc38),
		.ret_ras_index(DUT_ret_ras_index),

	    // update control
		.update_valid(tb_update_valid),
		.update_ras_index(tb_update_ras_index)
	);

    // ----------------------------------------------------------------
    // tasks:

    task check_outputs();
    begin
		if (expected_ret_pc38 !== DUT_ret_pc38) begin
			$display("TB ERROR: expected_ret_pc38 (%h) != DUT_ret_pc38 (%h)",
				expected_ret_pc38, DUT_ret_pc38);
			num_errors++;
			tb_error = 1'b1;
		end

		if (expected_ret_ras_index !== DUT_ret_ras_index) begin
			$display("TB ERROR: expected_ret_ras_index (%h) != DUT_ret_ras_index (%h)",
				expected_ret_ras_index, DUT_ret_ras_index);
			num_errors++;
			tb_error = 1'b1;
		end

        #(PERIOD / 10);
        tb_error = 1'b0;
    end
    endtask

    // ----------------------------------------------------------------
    // initial block:

    initial begin

        // ------------------------------------------------------------
        // reset:
        test_case = "reset";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

        // inputs:
        sub_test_case = "assert reset";
        $display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b0;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b0;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(posedge CLK); #(PERIOD/10);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h0000000000;
		expected_ret_ras_index = 4'h0;
	    // update control

		check_outputs();

        // inputs:
        sub_test_case = "deassert reset";
        $display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b0;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(posedge CLK); #(PERIOD/10);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h0000000000;
		expected_ret_ras_index = 4'h0;
	    // update control

		check_outputs();

        // ------------------------------------------------------------
        // simple chain:
        test_case = "simple chain";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "link 1";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b1;
		tb_link_pc38 = 38'h1111111111;
	    // pc_gen return control
		tb_ret_valid = 1'b0;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h0000000000;
		expected_ret_ras_index = 4'h0;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "link 2";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // RESP stage
	    // pc_gen link control
		tb_link_valid = 1'b1;
		tb_link_pc38 = 38'h2222222222;
	    // pc_gen return control
		tb_ret_valid = 1'b0;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h1111111111;
		expected_ret_ras_index = 4'h1;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "ret 2";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h3333333333;
	    // pc_gen return control
		tb_ret_valid = 1'b1;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h2222222222;
		expected_ret_ras_index = 4'h2;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "link + ret 1";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b1;
		tb_link_pc38 = 38'h5555555555;
	    // pc_gen return control
		tb_ret_valid = 1'b1;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h1111111111;
		expected_ret_ras_index = 4'h1;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "update to E";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b0;
	    // update control
		tb_update_valid = 1'b1;
		tb_update_ras_index = 4'hE;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h5555555555;
		expected_ret_ras_index = 4'h1;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "update to 3";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b0;
	    // update control
		tb_update_valid = 1'b1;
		tb_update_ras_index = 4'h3;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h0000000000;
		expected_ret_ras_index = 4'hE;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "ret to 2";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b1;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h0000000000;
		expected_ret_ras_index = 4'h3;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "ret to 1";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b1;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h2222222222;
		expected_ret_ras_index = 4'h2;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "ret to 0";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b1;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h5555555555;
		expected_ret_ras_index = 4'h1;
	    // update control

		check_outputs();

		@(posedge CLK); #(PERIOD/10);

		// inputs
		sub_test_case = "done";
		$display("\t- sub_test: %s", sub_test_case);

		// reset
		nRST = 1'b1;
	    // pc_gen link control
		tb_link_valid = 1'b0;
		tb_link_pc38 = 38'h0000000000;
	    // pc_gen return control
		tb_ret_valid = 1'b0;
	    // update control
		tb_update_valid = 1'b0;
		tb_update_ras_index = 4'h0;

		@(negedge CLK);

		// outputs:

	    // pc_gen link control
	    // pc_gen return control
		expected_ret_pc38 = 38'h0000000000;
		expected_ret_ras_index = 4'h0;
	    // update control

		check_outputs();

        // ------------------------------------------------------------
        // finish:
        @(posedge CLK); #(PERIOD/10);
        
        test_case = "finish";
        $display("\ntest %0d: %s", test_num, test_case);
        test_num++;

        @(posedge CLK); #(PERIOD/10);

        $display();
        if (num_errors) begin
            $display("FAIL: %d tests fail", num_errors);
        end
        else begin
            $display("SUCCESS: all tests pass");
        end
        $display();

        $finish();
    end

endmodule