module alu_reg_mdu_iq_sva ();
    
endmodule